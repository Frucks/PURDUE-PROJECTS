// $Id: $
// File name:   tb_flex_counter.sv
// Created:     2/1/2023
// Author:      Joao Taff-Freire
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: .

// 0.5um D-FlipFlop Timing Data Estimates:
// Data Propagation delay (clk->Q): 670ps
// Setup time for data relative to clock: 190ps
// Hold time for data relative to clock: 10ps

`timescale 10ns / 100ps

module tb_flex_counter();

  // Define local parameters used by the test bench
  localparam  CLK_PERIOD    = 1;
  localparam  FF_SETUP_TIME = 0.190;
  localparam  FF_HOLD_TIME  = 0.100;
  localparam  CHECK_DELAY   = (CLK_PERIOD - FF_SETUP_TIME); // Check right before the setup time starts
  
  localparam  INACTIVE_VALUE     = '0;
  localparam  RESET_OUTPUT_VALUE = INACTIVE_VALUE;

  localparam NUM_CNT_BIT = 4;
  
  // Declare DUT portmap signals
  reg tb_clk;
  reg tb_n_rst;
  reg tb_clear;
  reg tb_count_enable;
  reg [NUM_CNT_BIT - 1:0] tb_rollover_val;
  wire [NUM_CNT_BIT - 1:0] tb_count_out;
  wire tb_rollover_flag;
  
  // Declare test bench signals
  integer tb_test_num;
  string tb_test_case;
  integer tb_stream_test_num;
  string tb_stream_check_tag;
  
  // Task for standard DUT reset procedure
  task reset_dut;
  begin
    // Activate the reset
    tb_n_rst = 1'b0;

    // Maintain the reset for more than one cycle
    @(posedge tb_clk);
    @(posedge tb_clk);

    // Wait until safely away from rising edge of the clock before releasing
    @(negedge tb_clk);
    tb_n_rst = 1'b1;

    // Leave out of reset for a couple cycles before allowing other stimulus
    // Wait for negative clock edges, 
    // since inputs to DUT should normally be applied away from rising clock edges
    @(negedge tb_clk);
    @(negedge tb_clk);
  end
  endtask

  task clear_dut;
  begin
    // Activate the clear
    @(negedge tb_clk);
    tb_clear = 1'b1;

    // Maintain the clear for one cycle
    @(posedge tb_clk);

    // Wait until safely away from rising edge of the clock before releasing
    @(negedge tb_clk);
    tb_clear = 1'b0;
  end
  endtask

  // Task to cleanly and consistently check DUT output values
  task check_output;
    input logic  [NUM_CNT_BIT - 1:0] expected_value;
    input string check_tag;
  begin
    if(expected_value == tb_count_out) begin // Check passed
      $info("Correct counter output %s during %s test case", check_tag, tb_test_case);
    end
    else begin // Check failed
      $error("Incorrect counter output %s during %s test case", check_tag, tb_test_case);
    end
  end
  endtask

  task check_flag;
   input logic  expected_value;
   input string check_tag;
  begin
    if(expected_value == tb_rollover_flag) begin // Check passed
      $info("Correct rollover flag %s during %s test case", check_tag, tb_test_case);
    end
    else begin // Check failed
      $error("Incorrect rollover flag %s during %s test case", check_tag, tb_test_case);
    end
  end
  endtask

//   // Task to cleanly and consistently check for correct values during MetaStability Test Cases
//   task check_output_meta;
//     input string check_tag;
//   begin
//     // Only need to check that it's not a metastable value since decays are random
//     if((1'b1 == tb_sync_out) || (1'b0 == tb_sync_out)) begin // Check passed
//       $info("Correct synchronizer output %s during %s test case", check_tag, tb_test_case);
//     end
//     else begin // Check failed
//       $error("Incorrect synchronizer output %s during %s test case", check_tag, tb_test_case);
//     end
//   end
//   endtask

  // Clock generation block
  always
  begin
    // Start with clock low to avoid false rising edge events at t=0
    tb_clk = 1'b0;
    // Wait half of the clock period before toggling clock value (maintain 50% duty cycle)
    #(CLK_PERIOD/2.0);
    tb_clk = 1'b1;
    // Wait half of the clock period before toggling clock value via rerunning the block (maintain 50% duty cycle)
    #(CLK_PERIOD/2.0);
  end
  
  // DUT Port map
  flex_counter DUT (.clk(tb_clk), .n_rst(tb_n_rst), .clear(tb_clear), .count_enable(tb_count_enable), .rollover_val(tb_rollover_val), .count_out(tb_count_out), .rollover_flag(tb_rollover_flag));
  
  // Test bench main process
  initial
  begin
    // Initialize all of the test inputs
    tb_n_rst  = 1'b1;              // Initialize to be inactive
    tb_count_enable  = INACTIVE_VALUE; // Initialize input to inactive  value
    tb_test_num = 0;               // Initialize test case counter
    tb_test_case = "Test bench initializaton";
    tb_stream_test_num = 0;
    tb_stream_check_tag = "N/A";
    tb_clear = 'd0;
    tb_rollover_val = 'd0;
    // Wait some time before starting first test case
    #(0.1);
    
    // ************************************************************************
    // Test Case 1: Power-on Reset of the DUT
    // ************************************************************************
    tb_test_num = tb_test_num + 1;
    tb_test_case = "Power on Reset";
    // Note: Do not use reset task during reset test case since we need to specifically check behavior during reset
    // Wait some time before applying test case stimulus
    #(0.1);
    // Apply test case initial stimulus
    tb_count_enable  = INACTIVE_VALUE; // Set to be the the non-reset value
    tb_n_rst  = 1'b0;    // Activate reset
    
    // Wait for a bit before checking for correct functionality
    #(CLK_PERIOD * 0.5);

    // Check that internal state was correctly reset
    check_output( RESET_OUTPUT_VALUE, 
                  "after reset applied");
    
    // Check that the reset value is maintained during a clock cycle
    #(CLK_PERIOD);
    check_output( RESET_OUTPUT_VALUE, 
                  "after clock cycle while in reset");
    
    // Release the reset away from a clock edge
    @(posedge tb_clk);
    #(2 * FF_HOLD_TIME);
    tb_n_rst  = 1'b1;   // Deactivate the chip reset
    #0.1;
    // Check that internal state was correctly keep after reset release
    check_output( RESET_OUTPUT_VALUE, 
                  "after reset was released");

    // ************************************************************************    
    // Test Case 2: Rollover for a rollover value that is not a power of two
    // ************************************************************************
    @(negedge tb_clk); 
    tb_test_num = tb_test_num + 1;
    tb_test_case = "Rollover for a rollover value that is not a power of two";
    // Start out with inactive value and reset the DUT to isolate from prior tests
    tb_count_enable = INACTIVE_VALUE;
    reset_dut();

    // Assign test case stimulus
    tb_rollover_val = 'd3;
    tb_count_enable = 1'b1;

    // Wait for DUT to process stimulus before checking results
    @(posedge tb_clk); 
    @(posedge tb_clk); 
    @(posedge tb_clk);
    #(CHECK_DELAY);
    check_output( tb_rollover_val,
                  "after processing delay");
    check_flag( 1'b1,
                  "after processing delay");
    @(posedge tb_clk); 
    // Move away from risign edge and allow for propagation delays before checking
    #(CHECK_DELAY);
    // Check results
    check_output( 1'b1,
                  "after processing delay");
    check_flag( 1'b0,
                  "after processing delay");
    
    // ************************************************************************    
    // Test Case 3: Continuous counting
    // ************************************************************************
    @(negedge tb_clk); 
    tb_test_num = tb_test_num + 1;
    tb_test_case = "Continuous counting";
    // Start out with inactive value and reset the DUT to isolate from prior tests
    tb_count_enable = INACTIVE_VALUE;
    reset_dut();

    // Assign test case stimulus
    tb_rollover_val = 2 ** (NUM_CNT_BIT) - 1;
    tb_count_enable = 1'b1;

    // Wait for DUT to process stimulus before checking results
    for (int i = 1; i < tb_rollover_val; i++) begin
      #(CHECK_DELAY);
      check_output( i,
                "after processing delay");
       check_flag( 1'b0,
                "afterprocessing delay");
      @(posedge tb_clk);
    end
    #(CHECK_DELAY);
    check_output( tb_rollover_val,
                  "after processing delay");
    check_flag( 1'b1,
                  "after processing delay");
    @(posedge tb_clk);
    #(CHECK_DELAY);
    check_output( 'd1,
                  "after processing delay");
    check_flag( 1'b0,
                  "after processing delay");
    
    // ************************************************************************    
    // Test Case 4: Discontinuous counting
    // ************************************************************************
      @(negedge tb_clk); 
    tb_test_num = tb_test_num + 1;
    tb_test_case = "Discontinuous counting";
    // Start out with inactive value and reset the DUT to isolate from prior tests
    tb_count_enable = INACTIVE_VALUE;
    reset_dut();

    // Assign test case stimulus
    tb_rollover_val = 'd3;
    tb_count_enable = 1'b1;

    // Wait for DUT to process stimulus before checking results
    @(posedge tb_clk);
    #(CHECK_DELAY);
    check_output( 'd1,
                  "after processing delay");
    check_flag( 1'b0,
                  "after processing delay");
    @(posedge tb_clk);
    #(CHECK_DELAY);
    check_output( 'd2,
                  "after processing delay");
    check_flag( 1'b0,
                  "after processing delay");
    @(posedge tb_clk);
    #(CHECK_DELAY);
    check_output( 'd3,
                  "after processing delay");
    check_flag( 1'b1,
                  "after processing delay");
    tb_count_enable = 1'b0;
    @(posedge tb_clk);
    #(CHECK_DELAY);
    check_output( 'd3,
                  "after processing delay");
    check_flag( 1'b1,
                  "after processing delay");
    tb_count_enable = 1'b1;
    @(posedge tb_clk);
    #(CHECK_DELAY);
    check_output( 'd1,
                  "after processing delay");
    check_flag( 1'b0,
                  "after processing delay");

    // ************************************************************************    
    // Test Case 5: Clearing while counting to check clear vs. count enable priority
    // ************************************************************************
    @(negedge tb_clk); 
    tb_test_num = tb_test_num + 1;
    tb_test_case = "Clearing while counting";
    // Start out with inactive value and reset the DUT to isolate from prior tests
    tb_count_enable = INACTIVE_VALUE;
    reset_dut();

    // Assign test case stimulus
    tb_rollover_val = 'd3;
    tb_count_enable = 1'b1;

    // Wait for DUT to process stimulus before checking results
    @(posedge tb_clk);
    @(posedge tb_clk);
    clear_dut();
    @(posedge tb_clk);
    #(CHECK_DELAY);
    check_output( 'd1,
                  "after processing delay");
    check_flag( 1'b0,
                  "after processing delay");
    @(posedge tb_clk);
    #(CHECK_DELAY);
    check_output( 'd2,
                  "after processing delay");
    check_flag( 1'b0,
                  "after processing delay");
    $stop;   
  end
endmodule